// dj_tb.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module dj_tb (
	);

	wire         dj_inst_sc_fifo_0_almost_empty_data; // dj_inst:sc_fifo_0_almost_empty_data -> dj_inst_sc_fifo_0_almost_empty_bfm:sink_data
	wire         dj_inst_sc_fifo_0_almost_full_data;  // dj_inst:sc_fifo_0_almost_full_data -> dj_inst_sc_fifo_0_almost_full_bfm:sink_data
	wire         dj_inst_sc_fifo_0_out_valid;         // dj_inst:sc_fifo_0_out_valid -> dj_inst_sc_fifo_0_out_bfm:sink_valid
	wire  [15:0] dj_inst_sc_fifo_0_out_data;          // dj_inst:sc_fifo_0_out_data -> dj_inst_sc_fifo_0_out_bfm:sink_data
	wire         dj_inst_sc_fifo_0_out_ready;         // dj_inst_sc_fifo_0_out_bfm:sink_ready -> dj_inst:sc_fifo_0_out_ready
	wire   [0:0] dj_inst_sc_fifo_0_in_bfm_src_valid;  // dj_inst_sc_fifo_0_in_bfm:src_valid -> dj_inst:sc_fifo_0_in_valid
	wire  [15:0] dj_inst_sc_fifo_0_in_bfm_src_data;   // dj_inst_sc_fifo_0_in_bfm:src_data -> dj_inst:sc_fifo_0_in_data
	wire         dj_inst_sc_fifo_0_in_bfm_src_ready;  // dj_inst:sc_fifo_0_in_ready -> dj_inst_sc_fifo_0_in_bfm:src_ready
	wire         dj_inst_clk_bfm_clk_clk;             // dj_inst_clk_bfm:clk -> [dj_inst:clk_clk, dj_inst_reset_bfm:clk, dj_inst_sc_fifo_0_almost_empty_bfm:clk, dj_inst_sc_fifo_0_almost_full_bfm:clk, dj_inst_sc_fifo_0_in_bfm:clk, dj_inst_sc_fifo_0_out_bfm:clk]
	wire         dj_inst_reset_bfm_reset_reset;       // dj_inst_reset_bfm:reset -> [dj_inst:reset_reset_n, dj_inst_sc_fifo_0_almost_empty_bfm:reset, dj_inst_sc_fifo_0_almost_full_bfm:reset, dj_inst_sc_fifo_0_in_bfm:reset, dj_inst_sc_fifo_0_out_bfm:reset]

	dj dj_inst (
		.clk_clk                     (dj_inst_clk_bfm_clk_clk),             //                    clk.clk
		.reset_reset_n               (dj_inst_reset_bfm_reset_reset),       //                  reset.reset_n
		.sc_fifo_0_almost_empty_data (dj_inst_sc_fifo_0_almost_empty_data), // sc_fifo_0_almost_empty.data
		.sc_fifo_0_almost_full_data  (dj_inst_sc_fifo_0_almost_full_data),  //  sc_fifo_0_almost_full.data
		.sc_fifo_0_in_data           (dj_inst_sc_fifo_0_in_bfm_src_data),   //           sc_fifo_0_in.data
		.sc_fifo_0_in_valid          (dj_inst_sc_fifo_0_in_bfm_src_valid),  //                       .valid
		.sc_fifo_0_in_ready          (dj_inst_sc_fifo_0_in_bfm_src_ready),  //                       .ready
		.sc_fifo_0_out_data          (dj_inst_sc_fifo_0_out_data),          //          sc_fifo_0_out.data
		.sc_fifo_0_out_valid         (dj_inst_sc_fifo_0_out_valid),         //                       .valid
		.sc_fifo_0_out_ready         (dj_inst_sc_fifo_0_out_ready)          //                       .ready
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dj_inst_clk_bfm (
		.clk (dj_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dj_inst_reset_bfm (
		.reset (dj_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dj_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (0),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (0),
		.USE_VALID        (0),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (1),
		.ST_NUMSYMBOLS    (1),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (1),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) dj_inst_sc_fifo_0_almost_empty_bfm (
		.clk                (dj_inst_clk_bfm_clk_clk),             //       clk.clk
		.reset              (~dj_inst_reset_bfm_reset_reset),      // clk_reset.reset
		.sink_data          (dj_inst_sc_fifo_0_almost_empty_data), //      sink.data
		.sink_valid         (1'b1),                                // (terminated)
		.sink_ready         (),                                    // (terminated)
		.sink_startofpacket (1'b0),                                // (terminated)
		.sink_endofpacket   (1'b0),                                // (terminated)
		.sink_empty         (1'b0),                                // (terminated)
		.sink_channel       (1'b0),                                // (terminated)
		.sink_error         (1'b0)                                 // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (0),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (0),
		.USE_VALID        (0),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (1),
		.ST_NUMSYMBOLS    (1),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (1),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (1)
	) dj_inst_sc_fifo_0_almost_full_bfm (
		.clk                (dj_inst_clk_bfm_clk_clk),            //       clk.clk
		.reset              (~dj_inst_reset_bfm_reset_reset),     // clk_reset.reset
		.sink_data          (dj_inst_sc_fifo_0_almost_full_data), //      sink.data
		.sink_valid         (1'b1),                               // (terminated)
		.sink_ready         (),                                   // (terminated)
		.sink_startofpacket (1'b0),                               // (terminated)
		.sink_endofpacket   (1'b0),                               // (terminated)
		.sink_empty         (1'b0),                               // (terminated)
		.sink_channel       (1'b0),                               // (terminated)
		.sink_error         (1'b0)                                // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (0),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (2),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (1),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) dj_inst_sc_fifo_0_in_bfm (
		.clk               (dj_inst_clk_bfm_clk_clk),            //       clk.clk
		.reset             (~dj_inst_reset_bfm_reset_reset),     // clk_reset.reset
		.src_data          (dj_inst_sc_fifo_0_in_bfm_src_data),  //       src.data
		.src_valid         (dj_inst_sc_fifo_0_in_bfm_src_valid), //          .valid
		.src_ready         (dj_inst_sc_fifo_0_in_bfm_src_ready), //          .ready
		.src_startofpacket (),                                   // (terminated)
		.src_endofpacket   (),                                   // (terminated)
		.src_empty         (),                                   // (terminated)
		.src_channel       (),                                   // (terminated)
		.src_error         ()                                    // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (0),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (2),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (1),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (2)
	) dj_inst_sc_fifo_0_out_bfm (
		.clk                (dj_inst_clk_bfm_clk_clk),        //       clk.clk
		.reset              (~dj_inst_reset_bfm_reset_reset), // clk_reset.reset
		.sink_data          (dj_inst_sc_fifo_0_out_data),     //      sink.data
		.sink_valid         (dj_inst_sc_fifo_0_out_valid),    //          .valid
		.sink_ready         (dj_inst_sc_fifo_0_out_ready),    //          .ready
		.sink_startofpacket (1'b0),                           // (terminated)
		.sink_endofpacket   (1'b0),                           // (terminated)
		.sink_empty         (1'b0),                           // (terminated)
		.sink_channel       (1'b0),                           // (terminated)
		.sink_error         (1'b0)                            // (terminated)
	);


	always begin
		#10 clk <= ~clk;
	end

	initial begin
		dj_inst_clk_bfm_clk_clk <= 1'b0;
		dj_inst_clk_bfm_reset_reset <= 1'b1;
		#30 dj_inst_clk_bfm_reset_reset <= 1'b0;
		
	end

endmodule
